module approx_multiplier();
   



endmodule: approx_multiplier
